`include "Memory/Memory Module/memory.v"

module memory_tb;

endmodule