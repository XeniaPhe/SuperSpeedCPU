`timescale 1ns/1ns
`include "Control Unit/Control Unit/control_unit.v"

module control_unit_tb;
    
endmodule