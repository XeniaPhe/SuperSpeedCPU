`include "Control Unit/Instruction Decoder/instruction_decoder.v"

module instruction_decoder_tb;

endmodule