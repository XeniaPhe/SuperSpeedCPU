`include "Latches/Rising Edge Triggered D Flip-Flop/rising_edge_triggered_d_flipflop.v"
`include "Latches/Falling Edge Triggered D Flip-Flop/falling_edge_triggered_d_flipflop.v"

module terminator(
    input decode, halt_instruction, stack_overflow, instruction_end, pc_overflow, clk,
    output halted);

    

endmodule